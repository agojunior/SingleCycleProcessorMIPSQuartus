module  Instructions (PC,Inst, clock);

input clock;
output   [31:0] Inst;
input 	[10:0] PC;
reg 		[31:0] ramInstrucoes [31:0];
//always @(posedge clock) begin
initial begin
	//IN OUT DEMONSTRATION
	//ramInstrucoes[0] = 32'b01100000000000010000000000000110; //li r1, 6
	//ramInstrucoes[1] = {{6'b001110},{5'b00000},{5'b00011},{5'b00000},{5'b00000},{6'b000000}}; //in r3
	//ramInstrucoes[2] = {{6'b001111},{5'b00000},{5'b00001},{5'b00000},{5'b00000},{6'b000000}}; //out r1
	//ramInstrucoes[3] = {{6'b001111},{5'b00000},{5'b00011},{5'b00000},{5'b00000},{6'b000000}}; //out r3
	//ramInstrucoes[4] = {{6'b010000},{5'b00000},{5'b00000},{5'b00000},{5'b00000},{6'b000001}}; //j 1
	
	//ramInstrucoes[3] = 32'b00000000010000100001000000000111; //shl r2, r2, r2
	//ramInstrucoes[4] = {{6'b000000},{5'b00001},{5'b00010},{5'b00001},{5'b00000},{6'b000001}}; //sub r1, r2, r1
	//ramInstrucoes[5] = {{6'b000000},{5'b00010},{5'b00001},{5'b00011},{5'b00000},{6'b000001}}; //sub r2, r1, r3
	//ramInstrucoes[6] = {{6'b001101},{5'b00000},{5'b00010},{5'b00000},{5'b00000},{6'b000010}}; //sr r2, 2
	//ramInstrucoes[7] = {{6'b001100},{5'b00000},{5'b00010},{5'b00000},{5'b00000},{6'b000010}}; //lr r2, 2
	//ramInstrucoes[8] = {{6'b010000},{5'b00000},{5'b00000},{5'b00000},{5'b00000},{6'b000010}}; //j 2
	
	//FIBONACCI
	//ramInstrucoes[0] = {{6'b001110},{5'b00000},{5'b00001},{5'b00000},{5'b00000},{6'b000000}}; //in r3
	//FIBONACCI
	ramInstrucoes[0] = {{6'b001110},{5'b00000},{5'b00100},{5'b00000},{5'b00000},{6'b000000}}; //in r4
	//ramInstrucoes[0] = {{6'b011000},{5'b00000},{5'b00100},{5'b00000},{5'b00000},{6'b000101}}; //li r4,5
	ramInstrucoes[1] = {{6'b011000},{5'b00000},{5'b00001},{5'b00000},{5'b00000},{6'b000000}}; //li r1,0
	ramInstrucoes[2] = {{6'b011000},{5'b00000},{5'b00010},{5'b00000},{5'b00000},{6'b000001}}; //li r2,1
	ramInstrucoes[3] = {{6'b011000},{5'b00000},{5'b00101},{5'b00000},{5'b00000},{6'b000001}}; //li r5,1
	ramInstrucoes[4] = {{6'b000000},{5'b00010},{5'b00001},{5'b00011},{5'b00000},{6'b000000}}; //add  r1, r2, r3
	ramInstrucoes[5] = {{6'b001000},{5'b00010},{5'b00001},{5'b00000},{5'b00000},{6'b000000}}; //addi r2, rd1, 0
	ramInstrucoes[6] = {{6'b001001},{5'b00011},{5'b00010},{5'b00000},{5'b00000},{6'b000000}}; //subi r3,rd2,0
	ramInstrucoes[7] = {{6'b001000},{5'b00101},{5'b00101},{5'b00000},{5'b00000},{6'b000001}}; //addi r5, r5, 1
	ramInstrucoes[8] = {{6'b001010},{5'b00101},{5'b00100},{5'b00000},{5'b00000},{6'b000010}}; //beq r4,r5,2
	ramInstrucoes[9] = {{6'b001011},{5'b00101},{5'b00100},{16'b1111111111111011}}; //bnq r4,r5,-5
	ramInstrucoes[10] = {{6'b001111},{5'b00000},{5'b00011},{5'b00000},{5'b00000},{6'b000000}}; //out r3
	ramInstrucoes[11] = {{6'b111001},{5'b00001},{5'b00010},{5'b00011},{5'b00000},{6'b001010}}; //halt
end
assign Inst = ramInstrucoes[PC];

endmodule

//initial begin

	// $readmemb(".mif",ramInstrucoes);
	//end
